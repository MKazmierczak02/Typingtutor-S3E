library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_TEXTIO.ALL;

entity String_printer_2 is
    port ( Clk : in  STD_LOGIC;
           Reset : in  STD_LOGIC;
           TxBusy : in  STD_LOGIC;
           DIRdy : in  STD_LOGIC;              
           F0 : in  STD_LOGIC;
           DI : in STD_LOGIC_VECTOR (7 downto 0);
           DO : out  STD_LOGIC_VECTOR (7 downto 0);
           DORdy : out  STD_LOGIC;           
           Finished : out  STD_LOGIC;
           Busy : out  STD_LOGIC  );
end String_printer_2;

architecture RTL of String_printer_2 is

  -- FSM
  type state_type is (
    sReset,
    sBusyWait,
    sWE,
    sLoop,
    sReady,
    keyboardWait,
    sKeyboardWE,
    keyboardBusy,
    keyboardReady,
    keyboardFinished
    );
  signal State, nextState : state_type; 

  -- String to print
  type STRINGZ is array ( NATURAL range <> ) of CHARACTER;
  constant nStrSize : POSITIVE := 97;  
  constant textStrSize : POSITIVE := 49;

  signal romStr : STRINGZ( 0 to nStrSize - 1 ) := "Hello, it's typing tutor. Let's get it started! happy giraffe went to lorem ipsum dolor sit amet" & NUL;  
  signal keyboardStr : STRINGZ( 0 to textStrSize - 1 ) := "happy giraffe went to lorem ipsum dolor sit amet" & NUL;

  -- Character index
  signal cntIdx : std_logic_vector( 7 downto 0 ) := ( others => '0' );
  signal cntIdxKeyboard : std_logic_vector( 7 downto 0 ) := ( others => '0' );
  
  signal regDI : STD_LOGIC_VECTOR (7 downto 0);

begin
    
  regDI <= DI when rising_edge( Clk) and State = sReady;

  -- FSM
    process ( Clk )
    begin
        if rising_edge( Clk ) then
            if Reset = '1' then
                State <= sReset;
            else
                State <= nextState;
            end if;
            
            if State = sReset then
                cntIdxKeyboard <= ( others => '0' );
            elsif State = sWE then
                cntIdx <= cntIdx + 1;
            elsif State = sKeyboardWE then
                cntIdxKeyboard <= cntIdxKeyboard + 1;
            end if;
                        
        end if;
    end process;

    -- Function to map character to keycode
    function char_to_keycode(c : CHARACTER) return STD_LOGIC_VECTOR is
    begin
        case c is
            when 'A' => return "00011100";
            when 'B' => return "00110010";
            when 'C' => return "00100001";
            when 'D' => return "00100011";
            when 'E' => return "00100100";
            when 'F' => return "00101011";
            when 'G' => return "00110100";
            when 'H' => return "00110011";
            when 'I' => return "01000011";
            when 'J' => return "00111011";
            when 'K' => return "01000010";
            when 'L' => return "01001011";
            when 'M' => return "00111010";
            when 'N' => return "00110001";
            when 'O' => return "01000100";
            when 'P' => return "01001101";
            when 'Q' => return "00010101";
            when 'R' => return "00101101";
            when 'S' => return "00011011";
            when 'T' => return "00101100";
            when 'U' => return "00111100";
            when 'V' => return "00101010";
            when 'W' => return "00011101";
            when 'X' => return "00100010";
            when 'Y' => return "00110101";
            when 'Z' => return "00011010";
            when ' ' => return "00101001";
            when others => return "00000000"; -- Default for unsupported characters
        end case;
    end function;

    process( State, TxBusy, DIRdy, cntIdx, romStr, cntIdxKeyboard, keyboardStr, DI)
    begin
        nextState <= State;   -- default is to stay in current State
        
        case State is

            when sReset =>
                nextState <= sBusyWait;

            when sBusyWait =>
                if TxBusy = '0' then
                    nextState <= sWE;
                end if;

            when sWE =>   -- WE pulse
                nextState <= sLoop;

            when sReady =>
                if DIRdy = '1' then
                    nextState <= sWE;
                end if;
             
            when sLoop =>
                if romStr( conv_integer( cntIdx ) ) /= NUL then
                    nextState <= sBusyWait;
                else
                    nextState <= keyboardWait;
                end if;   

            when keyboardWait =>
                if DIRdy = '1' then
                    if DI = char_to_keycode(keyboardStr(conv_integer(cntIdxKeyboard))) then
                        if keyboardStr( conv_integer( cntIdxKeyboard ) ) /= NUL then
                            nextState <= keyboardReady;
                        else
                            nextState <= keyboardFinished;
                        end if;
                    end if;     
                end if;
                
            when keyboardReady =>
                if TxBusy = '0' then 
                    nextState <= sKeyboardWE;
                end if;
         
            when sKeyboardWE =>   -- WE pulse
                nextState <= keyboardBusy;
         
            when keyboardBusy =>
                if F0 = '0' then
                    nextState <= keyboardWait;
                end if;
                
            when keyboardFinished =>
                if F0 = '0' then
                    -- Handle finished state if needed
                end if;
            
        end case;
    end process;
          
    DORdy <= '1' when State = sWE OR State = sKeyboardWE else '0';  
    Finished <= '1' when State = keyboardFinished else '0';

    DO <= '0' & CONV_STD_LOGIC_VECTOR( CHARACTER'Pos( romStr( conv_integer( cntIdx ) ) ), 7 ) when (State = sBusyWait OR State = sWE OR State = sReady OR State = sLoop) else '0' & CONV_STD_LOGIC_VECTOR( CHARACTER'Pos( keyboardStr( conv_integer( cntIdxKeyboard ) ) ), 7 );
  
end RTL;
